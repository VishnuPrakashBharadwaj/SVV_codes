class generator;

endclass

