class receiver;

endclass

