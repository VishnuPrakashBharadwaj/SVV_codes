class scoreboard;

endclass

